
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Sbox8 is
port(

clk : in std_logic;
 rst : in std_logic;
 Sin: in std_logic_vector(5 downto 0);
 Sout : out std_logic_vector(3 downto 0) 


);



end Sbox8;

architecture Behavioral of Sbox8 is
signal temp : std_logic_vector(3 downto 0);
begin

process(clk,rst,Sin)

begin

 if rst='1' then
    temp<=(others=>'0');
   
 elsif clk'event and clk='1' then
     
	  case Sin is 
  -----------------------------------------------------------	  
  ----row #1 ------------------------------------------------
  -----------------------------------------------------------
        when "000000"=>
		     temp<="1101";
			  
			  
			when "000010"=>
           temp<="0010";			
			  
			  
			 when "000100"=>
            temp<="1000";			 
				
				
			 when "000110"=>
               temp<="0100";			 
					
					
			 when "001000"=>
               temp<="0110";			 
					
			 
			 when "001010"=>
                temp<="1111";			 
					 
					 
			  when "001100"=>
                temp<="1011";			  
					 
					 
			  when "001110"=>
                temp<="0001";			  
					 
				
            when "010000"=>
                 temp<="1010";				
					  
					  
				when "010010"=>
                  temp<="1001";				
						
						
				 when "010100"=>
                   temp<="0011";				 
						 
						 
				 when "010110"=>
                   temp<="1110";				 
						 
						 
				  when "011000"=>
                    temp<="0101";				  
						  
						  
					when "011010"=>
                    temp<="0000";					
						  
						
                when "011100"=>
                     temp<="1100";					 
							
							
					 when "011110"=>
                      temp<="0111";					 
							 
  -----------------------------------------------------------	  
  ----row #2 ------------------------------------------------
  -----------------------------------------------------------						 
				 
               when "000001"=>
                     temp<="0001";					
							
							
				    when "000011"=>
                      temp<="1111";					 
							 
							 
					  when "000101"=>
                       temp<="1101";					  
							  
							  
						when "000111"=>
                        temp<="1000";						
								
								
					    when "001001"=>
                         temp<="1010";						 
								 
								 
						  when "001011"=>
                          temp<="0011";						  
								  
								  
							when "001101"=>
                           temp<="0111";							
									
									
							when "001111"=>
                            temp<="0100";							 
  
                     
							when "010001"=>
                            temp<="1100";							
									 
									 
							when "010011"=>
                            temp<="0101";							
									 
									 
							when "010101"=>
                            temp<="0110";							
									 
									 
							when "010111"=>
                            temp<="1011";							
									 
									 
							when "011001"=>
                           temp<="0000";							
									
									
							 when "011011"=>
                           temp<="1110";							 
									
									
							  when "011101"=>
                            temp<="1001";							  
									 
									 
							  when "011111"=>
                             temp<="0010";							  
									  
  -----------------------------------------------------------	  
  ----row #3 ------------------------------------------------
  ----------
  -------------------------------------------------							  
	                   when "100000"=>
							       temp<="0111";
									 
							 when "100010"=>
                            temp<="1011";							 
									 
									 
							 when "100100"=>
                             temp<="0100";							 
									  
								
                       when "100110"=>
                             temp<="0001";							  
									  
									  
							  when "101000"=>
                              temp<="1001";							  
										
										
								when "101010"=>
                               temp<="1100";								
										 
										 
								 when "101100"=>
                                temp<="1110";								 
										  
										  
								 when "101110"=>
                                 temp<="0010";								 
											
								 when "110000"=>
                                  temp<="0000";								 
											 
								 when "110010"=>
                                   temp<="0110";								 
											  
											  
								 when "110100"=>
                                   temp<="1010";								 
											  
											  
								 when "110110"=>
                                    temp<="1101";								 
												
								  when "111000"=>
                                    temp<="1111";								  
												
												
									when "111010"=>
                                     temp<="0011";									
												 
												 
									when "111100"=>
                                      temp<="0101";									
												  
												  
									when "111110"=>
                                       temp<="1000";									
													
  -----------------------------------------------------------	  
  ----row #4 ------------------------------------------------
  -----------------------------------------------------------														
                            when "100001"=>
                                     temp<="0010";									 
												 
												 
									  when "100011"=>
                                     temp<="0001";									  
												 
												 
										when "100101"=>
                                     temp<="1110";										
												 
												 
										when "100111"=>
                                      temp<="0111";										


                               when "101001"=>
                                      temp<="0100";										 
												  
												  
										  when "101011"=>
                                      temp<="1010";										  
												  
												  
										  when "101101"=>
                                       temp<="1000";										  
													
													
										  when "101111"=>
                                       temp<="1101";										  
													
													
											when "110001"=>
                                       temp<="1111";											
													
													
											when "110011"=>
                                       temp<="1100"; 


                                 when "110101"=>
                                        temp<="1001";											
													 
													 
											when "110111"=>
                                         temp<="0000";											
													  
													  
											when "111001"=>
                                         temp<="0011";											
													  
											
                                  when "111011"=>
                                         temp<="0101";											 
													  
													  
											 when "111101"=>
                                          temp<="0110";											 
														
														
											 when "111111"=>
                                          temp<="1011";											 


          	
   -----------------------------------------------------------	  
  ----End of table-------------------------------------------
  -----------------------------------------------------------  			 
        when others =>		
		       temp <="0000";  
       
     end case;
  end if;	 
	 
	 

end process;



Sout<=temp;



















end Behavioral;

