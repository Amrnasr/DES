
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity PC1 is
port (

  
clk : in std_logic;

rst : in std_logic;

key : in std_logic_vector(63 downto 0);

PC1key : out std_logic_vector(55 downto 0) );



end PC1;

architecture Behavioral of PC1 is


signal temp : std_logic_vector(55 downto 0);

begin

process(clk,rst,key)
begin 

 if rst='1' then
 
   temp<=(others=>'0');
 
 elsif clk'event and clk='1' then
--  57 59 41 33 25 17 9
--	 1  58 50 42 34 26 18
--	 10 2  59 51 43 35 27
--	 19 11 3  60 52 44 36
--	 63 55 47 39 31 23 15
--	 7  62 54 46 38 30 22
--	 14 6  61 53 45 37 29
--	 21 13 5 28  20 12 4
 
 ------------------------------------------------
 --------------------first row in table-----------
 -------------------------------------------------
 temp(0)<=key(56);
 temp(1) <=key(58);
 temp(2) <= key(40);
 temp(3) <= key(32);
 temp(4) <= key(24);
 temp(5) <= key(16);
 temp(6) <= key(8);
 
 ----------------------------------------------------
 ----second row in table-------------------------------
 
 temp(7) <= key(0);
 temp(8) <= key(57);
 temp (9) <= key(49);
 temp(10) <= key(41);
 temp(11) <= key (33);
 temp(12) <=key(25);
 temp(13) <= key(26);
 
 -----------------------------------------------------
 --------------------------------------------third row
 -----------------------------------------------------
 --	 10 2  59 51 43 35 27
 
 temp(14) <=key(9);
 temp(15) <= key(1);
 temp(16) <= key(58);
 temp(17) <= key(50);
 temp(18) <= key(42);
 temp(19) <= key(34);
 temp(20) <= key(26);
 
 ---------------------------------------------------------
 ------------------------------------------------------
 -------------fourth row --------------------------------
 ---------------------------------------------------------
 ---------------------------------------------------------
 --	 19 11 3  60 52 44 36
 
 temp(21) <=key(18);
 temp(22) <= key(10);
 temp(23) <=key(2);
 temp(24) <= key(59);
 temp(25) <= key(51);
 temp(26) <= key(43);
 temp(27) <= key(35);
 --------------------------------------------------------
 ----------------------------------------------------------
 ---------------------------------------------------------
 -------fifth row-----------------------------------------
 ---------------------------------------------------------
 --	 63 55 47 39 31 23 15
 
 temp(28) <= key(62);
 temp(29) <= key(54);
 temp(30) <= key(46);
 temp(31) <= key(38);
 temp(32) <= key(30);
 temp(33) <= key(22);
 temp(34) <= key(14);
 
 ------------------------------------------------------------
 ------------------------------------------------------------
 -------------------------------------------------------------
 ----sixth row-----------------------------------------------
 -----------------------------------------------------------
 --	 7  62 54 46 38 30 22
 
 temp(35) <= key(6);
 temp(36) <= key(61);
 temp(37) <= key(53);
 temp(38) <= key(45);
 temp(39) <= key(37);
 temp(40) <= key(29);
 temp(41) <= key(21);
 
 --------------------------------------------------------------
 ------------------seventh row---------------------------------
 --------------------------------------------------------------
 --	 14 6  61 53 45 37 29

temp(42) <= key(13);
temp(43) <= key(5);
temp(44) <= key(60);
temp(45) <= key(52);
temp(46) <= key (44);
temp(47) <= key (36);
temp(48) <= key(28);


----------------------------------------------------
----------------------------------------------------
----------eighth row ------------------------------
---------------------------------------------------
---------------------------------------------------
--	 21 13 5 28  20 12 4----------------------------

temp(49) <= key(20);
temp(50) <= key(12);
temp(51) <= key(4);
temp(52) <= key(27);
temp(53) <= key(19);
temp(54) <= key(11);
temp(55) <=key(3);
 
 
 
 
 
 
 end if;




end process;


PC1key <=temp;

end Behavioral;

