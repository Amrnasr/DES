
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


entity IP-1 is
    Port ( clk : in  STD_LOGIC;
           input : in  STD_LOGIC_VECTOR (63 downto 0);
           output : out  STD_LOGIC_VECTOR (63 downto 0));
end IP-1;

architecture Behavioral of IP-1 is

begin







end Behavioral;

