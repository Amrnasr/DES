
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity PC2 is
port (

  
clk : in std_logic;

rst : in std_logic;

key : in std_logic_vector(55 downto 0);

PC2key : out std_logic_vector(47 downto 0) );


end PC2;

architecture Behavioral of PC2 is
signal temp : std_logic_vector(47 downto 0);
begin

process(clk,rst,key)

begin


--14 17 11 24 1  5  3 28 
--15 6 21  10 23 19 12 4
--26 8 16  7  27 20 13 2
--41 52 31 37 47 55 30 40
--51 45 33 48 44 49 39 56
--34 53 46 42 50 36 29 32


if rst='1' then


 temp<=(others=>'0');

elsif clk'event and clk='1' then
  --14 17 11 24 1  5  3 28 --------------
  ---row #1 -----------------------------
  ---------------------------------------
  
  temp(0) <= key(13);
  temp(1) <= key(16);
  temp(2) <= key(10);
  temp(3) <= key(23);
  temp(4) <= key(0);
  temp(5) <= key(4);
  temp(6) <= key(2);
  temp(7) <= key(27);
  
--15 6 21  10 23 19 12 4-----------------
----row #2 ------------------------------
temp(8) <= key(14);
temp(9) <= key(5);
temp(10) <=key(20);
temp(11) <=key(9);
temp(12) <=key(22);
temp(13) <=key(18);
temp(14) <=key(11);
temp(15) <=key(3);

-------------------------------------------------
-------------------------------------------------
-------------------------------------------------
--26 8 16  7  27 20 13 2-------------------------
----row #3 --------------------------------------

temp(16) <= key(25);
temp(17) <= key(7);
temp(18) <= key(15);
temp(19) <= key(6);
temp(20) <= key(26);
temp(21) <= key(19);
temp(22) <= key(12);
temp(23) <= key(1);

----------------------------------------------------
----------------------------------------------------
-----------row #4 ----------------------------------
----------------------------------------------------
-----41 52 31 37 47 55 30 40------------------------


temp(24)<= key(40);
temp(25)<= key(51);
temp(26) <= key(30);
temp(27) <= key(36);
temp(28) <= key(46);
temp(29) <= key(54);
temp(30) <= key(29);
temp(31) <= key(39);

----row #5------------------------------------------
--51 45 33 48 44 49 39 56---------------------------
----------------------------------------------------

temp(32) <= key(50);
temp(33) <= key(44);
temp(34) <= key(32);
temp(35) <= key(47);
temp(36) <= key(43);
temp(37) <= key(48);
temp(38) <= key(38);
temp(39) <= key(55);

---------------------------------------------------------
---------------------------------------------------------
---------------row #6 -----------------------------------
---------------------------------------------------------
--34 53 46 42 50 36 29 32

temp(40) <= key(33);
temp(41) <= key(52);
temp(42) <= key(45);
temp(43) <= key(41);
temp(44) <= key(49);
temp(45) <= key(35);
temp(46) <= key(28);
temp(47) <=key(31);
 
end if;

end process;

PC2key<=temp;

end Behavioral;

